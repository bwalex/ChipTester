module RingOscillator(output logic Q1,
                      input logic clock, Reset, Enable);

logic [3:0] count;

always_ff @(posedge clock, negedge Reset)
if(!Reset)
  begin
    Q1 = 0;
    count <= 0;
  end
else if(count == 4'b1000) count <=4'b0000;
else if(Enable)
  count <= count + 1;
else
  count <= 0;

always_ff @(posedge count[3], negedge Reset)
if(!Reset==0) Q1 <= 0;
else Q1 <= ~Q1;


endmodule