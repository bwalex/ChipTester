// sram_tb_bfm.v

// Generated using ACDS version 11.1sp2 259 at 2012.02.19.16:47:50

`timescale 1 ps / 1 ps
module sram_tb_bfm (
		output wire        sram_bridge_conduit_clock,       // sram_bridge_conduit.clock
		output wire [19:0] sram_bridge_conduit_address,     //                    .address
		output wire [1:0]  sram_bridge_conduit_byteenable,  //                    .byteenable
		input  wire [15:0] sram_bridge_conduit_readdata,    //                    .readdata
		output wire        sram_bridge_conduit_read,        //                    .read
		output wire        sram_bridge_conduit_write,       //                    .write
		output wire [15:0] sram_bridge_conduit_writedata,   //                    .writedata
		input  wire        sram_bridge_conduit_waitrequest  //                    .waitrequest
	);

	wire         reset_source_0_reset_reset;                                                                           // reset_source_0:reset -> [addr_router:reset, cmd_xbar_demux:reset, id_router:reset, mm_master_bfm_0:reset, mm_master_bfm_0_m0_translator:reset, mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:reset, rsp_xbar_demux:reset, sram_bridge_16_0:nreset, sram_bridge_16_0_avalon_slave_0_translator:reset, sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         clock_source_0_clk_clk;                                                                               // clock_source_0:clk -> [addr_router:clk, cmd_xbar_demux:clk, id_router:clk, mm_master_bfm_0:clk, mm_master_bfm_0_m0_translator:clk, mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:clk, reset_source_0:clk, rsp_xbar_demux:clk, sram_bridge_16_0:clock, sram_bridge_16_0_avalon_slave_0_translator:clk, sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire         mm_master_bfm_0_m0_waitrequest;                                                                       // mm_master_bfm_0_m0_translator:av_waitrequest -> mm_master_bfm_0:avm_waitrequest
	wire  [15:0] mm_master_bfm_0_m0_writedata;                                                                         // mm_master_bfm_0:avm_writedata -> mm_master_bfm_0_m0_translator:av_writedata
	wire  [19:0] mm_master_bfm_0_m0_address;                                                                           // mm_master_bfm_0:avm_address -> mm_master_bfm_0_m0_translator:av_address
	wire         mm_master_bfm_0_m0_write;                                                                             // mm_master_bfm_0:avm_write -> mm_master_bfm_0_m0_translator:av_write
	wire         mm_master_bfm_0_m0_read;                                                                              // mm_master_bfm_0:avm_read -> mm_master_bfm_0_m0_translator:av_read
	wire  [15:0] mm_master_bfm_0_m0_readdata;                                                                          // mm_master_bfm_0_m0_translator:av_readdata -> mm_master_bfm_0:avm_readdata
	wire   [1:0] mm_master_bfm_0_m0_byteenable;                                                                        // mm_master_bfm_0:avm_byteenable -> mm_master_bfm_0_m0_translator:av_byteenable
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest;                           // sram_bridge_16_0:waitrequest -> sram_bridge_16_0_avalon_slave_0_translator:av_waitrequest
	wire  [15:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                             // sram_bridge_16_0_avalon_slave_0_translator:av_writedata -> sram_bridge_16_0:writedata
	wire  [19:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                               // sram_bridge_16_0_avalon_slave_0_translator:av_address -> sram_bridge_16_0:address
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                 // sram_bridge_16_0_avalon_slave_0_translator:av_write -> sram_bridge_16_0:write
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_read;                                  // sram_bridge_16_0_avalon_slave_0_translator:av_read -> sram_bridge_16_0:read
	wire  [15:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                              // sram_bridge_16_0:readdata -> sram_bridge_16_0_avalon_slave_0_translator:av_readdata
	wire   [1:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;                            // sram_bridge_16_0_avalon_slave_0_translator:av_byteenable -> sram_bridge_16_0:byteenable
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // sram_bridge_16_0_avalon_slave_0_translator:uav_waitrequest -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;              // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_bridge_16_0_avalon_slave_0_translator:uav_burstcount
	wire  [15:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;               // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_bridge_16_0_avalon_slave_0_translator:uav_writedata
	wire  [20:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                 // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> sram_bridge_16_0_avalon_slave_0_translator:uav_address
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                   // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> sram_bridge_16_0_avalon_slave_0_translator:uav_write
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                    // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> sram_bridge_16_0_avalon_slave_0_translator:uav_lock
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                    // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> sram_bridge_16_0_avalon_slave_0_translator:uav_read
	wire  [15:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                // sram_bridge_16_0_avalon_slave_0_translator:uav_readdata -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // sram_bridge_16_0_avalon_slave_0_translator:uav_readdatavalid -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_bridge_16_0_avalon_slave_0_translator:uav_debugaccess
	wire   [1:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;              // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_bridge_16_0_avalon_slave_0_translator:uav_byteenable
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;            // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [52:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;             // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;            // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [52:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [15:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_waitrequest;                                  // mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> mm_master_bfm_0_m0_translator:uav_waitrequest
	wire   [1:0] mm_master_bfm_0_m0_translator_avalon_universal_master_0_burstcount;                                   // mm_master_bfm_0_m0_translator:uav_burstcount -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [15:0] mm_master_bfm_0_m0_translator_avalon_universal_master_0_writedata;                                    // mm_master_bfm_0_m0_translator:uav_writedata -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire  [20:0] mm_master_bfm_0_m0_translator_avalon_universal_master_0_address;                                      // mm_master_bfm_0_m0_translator:uav_address -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:av_address
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_lock;                                         // mm_master_bfm_0_m0_translator:uav_lock -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:av_lock
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_write;                                        // mm_master_bfm_0_m0_translator:uav_write -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:av_write
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_read;                                         // mm_master_bfm_0_m0_translator:uav_read -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:av_read
	wire  [15:0] mm_master_bfm_0_m0_translator_avalon_universal_master_0_readdata;                                     // mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:av_readdata -> mm_master_bfm_0_m0_translator:uav_readdata
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_debugaccess;                                  // mm_master_bfm_0_m0_translator:uav_debugaccess -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [1:0] mm_master_bfm_0_m0_translator_avalon_universal_master_0_byteenable;                                   // mm_master_bfm_0_m0_translator:uav_byteenable -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_readdatavalid;                                // mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> mm_master_bfm_0_m0_translator:uav_readdatavalid
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_valid;                               // mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [51:0] mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_data;                                // mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router:sink_ready -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                   // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [51:0] sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                    // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire         cmd_xbar_demux_src0_endofpacket;                                                                      // cmd_xbar_demux:src0_endofpacket -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                            // cmd_xbar_demux:src0_valid -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                    // cmd_xbar_demux:src0_startofpacket -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [51:0] cmd_xbar_demux_src0_data;                                                                             // cmd_xbar_demux:src0_data -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [0:0] cmd_xbar_demux_src0_channel;                                                                          // cmd_xbar_demux:src0_channel -> sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                      // rsp_xbar_demux:src0_endofpacket -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                            // rsp_xbar_demux:src0_valid -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                    // rsp_xbar_demux:src0_startofpacket -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [51:0] rsp_xbar_demux_src0_data;                                                                             // rsp_xbar_demux:src0_data -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:rp_data
	wire   [0:0] rsp_xbar_demux_src0_channel;                                                                          // rsp_xbar_demux:src0_channel -> mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire         addr_router_src_endofpacket;                                                                          // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                                // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                        // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [51:0] addr_router_src_data;                                                                                 // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [0:0] addr_router_src_channel;                                                                              // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                                // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_demux_src0_ready;                                                                            // mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src0_ready;                                                                            // sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire         id_router_src_endofpacket;                                                                            // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                  // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                          // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [51:0] id_router_src_data;                                                                                   // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [0:0] id_router_src_channel;                                                                                // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                  // rsp_xbar_demux:sink_ready -> id_router:src_ready

	altera_avalon_clock_source #(
		.CLOCK_RATE (100)
	) clock_source_0 (
		.clk (clock_source_0_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (1),
		.INITIAL_RESET_CYCLES (1)
	) reset_source_0 (
		.reset (reset_source_0_reset_reset), // reset.reset
		.clk   (clock_source_0_clk_clk)      //   clk.clk
	);

	altera_avalon_mm_master_bfm #(
		.AV_ADDRESS_W               (20),
		.AV_SYMBOL_W                (8),
		.AV_NUMSYMBOLS              (2),
		.AV_BURSTCOUNT_W            (1),
		.AV_READRESPONSE_W          (16),
		.AV_WRITERESPONSE_W         (16),
		.USE_READ                   (1),
		.USE_WRITE                  (1),
		.USE_ADDRESS                (1),
		.USE_BYTE_ENABLE            (1),
		.USE_BURSTCOUNT             (0),
		.USE_READ_DATA              (1),
		.USE_READ_DATA_VALID        (0),
		.USE_WRITE_DATA             (1),
		.USE_BEGIN_TRANSFER         (0),
		.USE_BEGIN_BURST_TRANSFER   (0),
		.USE_WAIT_REQUEST           (1),
		.USE_TRANSACTIONID          (0),
		.USE_WRITERESPONSE          (0),
		.USE_READRESPONSE           (0),
		.USE_CLKEN                  (0),
		.AV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_BURST_LINEWRAP          (1),
		.AV_BURST_BNDR_ONLY         (0),
		.AV_MAX_PENDING_READS       (0),
		.AV_FIX_READ_LATENCY        (0 /* was 1 */),
		.AV_READ_WAIT_TIME          (0 /* was 1 */),
		.AV_WRITE_WAIT_TIME         (0),
		.REGISTER_WAITREQUEST       (0),
		.AV_REGISTERINCOMINGSIGNALS (0)
	) mm_master_bfm_0 (
		.clk                      (clock_source_0_clk_clk),         //       clk.clk
		.reset                    (reset_source_0_reset_reset),     // clk_reset.reset
		.avm_address              (mm_master_bfm_0_m0_address),     //        m0.address
		.avm_readdata             (mm_master_bfm_0_m0_readdata),    //          .readdata
		.avm_writedata            (mm_master_bfm_0_m0_writedata),   //          .writedata
		.avm_waitrequest          (mm_master_bfm_0_m0_waitrequest), //          .waitrequest
		.avm_write                (mm_master_bfm_0_m0_write),       //          .write
		.avm_read                 (mm_master_bfm_0_m0_read),        //          .read
		.avm_byteenable           (mm_master_bfm_0_m0_byteenable),  //          .byteenable
		.avm_burstcount           (),                               // (terminated)
		.avm_begintransfer        (),                               // (terminated)
		.avm_beginbursttransfer   (),                               // (terminated)
		.avm_readdatavalid        (1'b0),                           // (terminated)
		.avm_arbiterlock          (),                               // (terminated)
		.avm_lock                 (),                               // (terminated)
		.avm_debugaccess          (),                               // (terminated)
		.avm_transactionid        (),                               // (terminated)
		.avm_readresponse         (16'b0000000000000000),           // (terminated)
		.avm_readid               (8'b00000000),                    // (terminated)
		.avm_writeresponserequest (),                               // (terminated)
		.avm_writeresponse        (16'b0000000000000000),           // (terminated)
		.avm_writeresponsevalid   (1'b0),                           // (terminated)
		.avm_writeid              (8'b00000000),                    // (terminated)
		.avm_clken                ()                                // (terminated)
	);

	sram_bridge #(
		.ADDR_WIDTH (20)
	) sram_bridge_16_0 (
		.byteenable    (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),  //           avalon_slave_0.byteenable
		.read          (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_read),        //                         .read
		.readdata      (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),    //                         .readdata
		.write         (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_write),       //                         .write
		.writedata     (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //                         .writedata
		.waitrequest   (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest), //                         .waitrequest
		.address       (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_address),     //                         .address
		.clock         (clock_source_0_clk_clk),                                                     //               clock_sink.clk
		.nreset        (~reset_source_0_reset_reset),                                                //               reset_sink.reset_n
		.m_clock       (sram_bridge_conduit_clock),                                                  // avalon_mm_master_conduit.export
		.m_address     (sram_bridge_conduit_address),                                                //                         .export
		.m_byteenable  (sram_bridge_conduit_byteenable),                                             //                         .export
		.m_readdata    (sram_bridge_conduit_readdata),                                               //                         .export
		.m_read        (sram_bridge_conduit_read),                                                   //                         .export
		.m_write       (sram_bridge_conduit_write),                                                  //                         .export
		.m_writedata   (sram_bridge_conduit_writedata),                                              //                         .export
		.m_waitrequest (sram_bridge_conduit_waitrequest)                                             //                         .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (20),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (21),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (0),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) mm_master_bfm_0_m0_translator (
		.clk                   (clock_source_0_clk_clk),                                                //                       clk.clk
		.reset                 (reset_source_0_reset_reset),                                            //                     reset.reset
		.uav_address           (mm_master_bfm_0_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (mm_master_bfm_0_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (mm_master_bfm_0_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (mm_master_bfm_0_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (mm_master_bfm_0_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (mm_master_bfm_0_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (mm_master_bfm_0_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (mm_master_bfm_0_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (mm_master_bfm_0_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (mm_master_bfm_0_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (mm_master_bfm_0_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (mm_master_bfm_0_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (mm_master_bfm_0_m0_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (mm_master_bfm_0_m0_byteenable),                                         //                          .byteenable
		.av_read               (mm_master_bfm_0_m0_read),                                               //                          .read
		.av_readdata           (mm_master_bfm_0_m0_readdata),                                           //                          .readdata
		.av_write              (mm_master_bfm_0_m0_write),                                              //                          .write
		.av_writedata          (mm_master_bfm_0_m0_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                  //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                  //               (terminated)
		.av_begintransfer      (1'b0),                                                                  //               (terminated)
		.av_chipselect         (1'b0),                                                                  //               (terminated)
		.av_readdatavalid      (),                                                                      //               (terminated)
		.av_lock               (1'b0),                                                                  //               (terminated)
		.av_debugaccess        (1'b0),                                                                  //               (terminated)
		.uav_clken             (),                                                                      //               (terminated)
		.av_clken              (1'b1)                                                                   //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (20),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sram_bridge_16_0_avalon_slave_0_translator (
		.clk                   (clock_source_0_clk_clk),                                                                     //                      clk.clk
		.reset                 (reset_source_0_reset_reset),                                                                 //                    reset.reset
		.uav_address           (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (sram_bridge_16_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_begintransfer      (),                                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                                           //              (terminated)
		.av_burstcount         (),                                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                                           //              (terminated)
		.av_lock               (),                                                                                           //              (terminated)
		.av_chipselect         (),                                                                                           //              (terminated)
		.av_clken              (),                                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                                       //              (terminated)
		.av_debugaccess        (),                                                                                           //              (terminated)
		.av_outputenable       ()                                                                                            //              (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (48),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (38),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (39),
		.PKT_TRANS_POSTED          (40),
		.PKT_TRANS_WRITE           (41),
		.PKT_TRANS_READ            (42),
		.PKT_TRANS_LOCK            (43),
		.PKT_SRC_ID_H              (49),
		.PKT_SRC_ID_L              (49),
		.PKT_DEST_ID_H             (50),
		.PKT_DEST_ID_L             (50),
		.PKT_BURSTWRAP_H           (47),
		.PKT_BURSTWRAP_L           (46),
		.PKT_BYTE_CNT_H            (45),
		.PKT_BYTE_CNT_L            (44),
		.PKT_PROTECTION_H          (51),
		.PKT_PROTECTION_L          (51),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (52),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clock_source_0_clk_clk),                                                                               //             clk.clk
		.reset                   (reset_source_0_reset_reset),                                                                           //       clk_reset.reset
		.m0_address              (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                                          //                .channel
		.rf_sink_ready           (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (53),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clock_source_0_clk_clk),                                                                               //       clk.clk
		.reset             (reset_source_0_reset_reset),                                                                           // clk_reset.reset
		.in_data           (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                                 // (terminated)
		.csr_readdata      (),                                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                 // (terminated)
		.almost_full_data  (),                                                                                                     // (terminated)
		.almost_empty_data (),                                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                                 // (terminated)
		.out_empty         (),                                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                                 // (terminated)
		.out_error         (),                                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                                 // (terminated)
		.out_channel       ()                                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (51),
		.PKT_PROTECTION_L          (51),
		.PKT_BEGIN_BURST           (48),
		.PKT_BURSTWRAP_H           (47),
		.PKT_BURSTWRAP_L           (46),
		.PKT_BYTE_CNT_H            (45),
		.PKT_BYTE_CNT_L            (44),
		.PKT_ADDR_H                (38),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (39),
		.PKT_TRANS_POSTED          (40),
		.PKT_TRANS_WRITE           (41),
		.PKT_TRANS_READ            (42),
		.PKT_TRANS_LOCK            (43),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (49),
		.PKT_SRC_ID_L              (49),
		.PKT_DEST_ID_H             (50),
		.PKT_DEST_ID_L             (50),
		.ST_DATA_W                 (52),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1)
	) mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent (
		.clk              (clock_source_0_clk_clk),                                                         //       clk.clk
		.reset            (reset_source_0_reset_reset),                                                     // clk_reset.reset
		.av_address       (mm_master_bfm_0_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (mm_master_bfm_0_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (mm_master_bfm_0_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (mm_master_bfm_0_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (mm_master_bfm_0_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (mm_master_bfm_0_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (mm_master_bfm_0_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (mm_master_bfm_0_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (mm_master_bfm_0_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (mm_master_bfm_0_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (mm_master_bfm_0_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_demux_src0_valid),                                                      //        rp.valid
		.rp_data          (rsp_xbar_demux_src0_data),                                                       //          .data
		.rp_channel       (rsp_xbar_demux_src0_channel),                                                    //          .channel
		.rp_startofpacket (rsp_xbar_demux_src0_startofpacket),                                              //          .startofpacket
		.rp_endofpacket   (rsp_xbar_demux_src0_endofpacket),                                                //          .endofpacket
		.rp_ready         (rsp_xbar_demux_src0_ready)                                                       //          .ready
	);

	sram_tb_bfm_addr_router addr_router (
		.sink_ready         (mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (mm_master_bfm_0_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clock_source_0_clk_clk),                                                         //       clk.clk
		.reset              (reset_source_0_reset_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_src_valid),                                                          //          .valid
		.src_data           (addr_router_src_data),                                                           //          .data
		.src_channel        (addr_router_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                     //          .endofpacket
	);

	sram_tb_bfm_id_router id_router (
		.sink_ready         (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_bridge_16_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clock_source_0_clk_clk),                                                                     //       clk.clk
		.reset              (reset_source_0_reset_reset),                                                                 // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                        //       src.ready
		.src_valid          (id_router_src_valid),                                                                        //          .valid
		.src_data           (id_router_src_data),                                                                         //          .data
		.src_channel        (id_router_src_channel),                                                                      //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                                //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                   //          .endofpacket
	);

	sram_tb_bfm_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clock_source_0_clk_clk),            //       clk.clk
		.reset              (reset_source_0_reset_reset),        // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	sram_tb_bfm_cmd_xbar_demux rsp_xbar_demux (
		.clk                (clock_source_0_clk_clk),            //       clk.clk
		.reset              (reset_source_0_reset_reset),        // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

endmodule
