module Inverter(output logic Q0,
                input logic A0);

assign Q0 = ~A0;

endmodule